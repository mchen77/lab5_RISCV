//intermediate generator module

module interm_gen();
endmodule
