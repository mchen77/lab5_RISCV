module lab05(clk, reset, foo);
	input clk;
	input reset;
	input foo;
	
	endmodule
	